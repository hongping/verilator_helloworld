module top();
  initial begin
    $display("hello world");
    $finish;
  end
endmodule : top